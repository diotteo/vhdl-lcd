----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:
-- Design Name:
-- Module Name:
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
use work.defs.all;

library IEEE;
use IEEE.std_logic_1164.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;



entity Set_Cgram_Address is
	port(
			clk : in std_logic;
			enable : in boolean;
			done : out boolean;
			address : in std_logic_vector(5 downto 0);
			lcd : out lcd_type
			);
end Set_Cgram_Address;


architecture Set_Cgram_Address of Set_Cgram_Address is
	signal instr : std_logic_vector(7 downto 0);
begin
	instr <= x"40" or address;

	COMP_WRITE : write_module port map (
			clk,
			enable,
			done,
			'0',
			instr,
			lcd
			);
end Set_Cgram_Address;
