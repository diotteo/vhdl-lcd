package defs is
	-- length in bits of the lcd vector
	constant LCD_LEN : integer := 11;
end package defs;

--package body defs is
--end package body defs;
