----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    10:15:18 01/27/2015
-- Design Name:
-- Module Name:    write_module - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;



entity write_module is
	port(
			clk : in    std_logic; --Signal de l'horloge cadenc� � 100Mhz

			-- Signaux permettant de contr�ler l'�tat du module
			send   : in  boolean; -- D�marre la s�quence d'envoie sur un front montant
			ins_in : in  std_logic_vector(8 downto 0); -- Instruction ou donn�e � envoyer(7 downto 0) + bit RS(8)
			done_write   : out boolean; -- Niveau haut lorsque le module a termin� l'envoie

			-- Signaux qui seront li�s au LCD
			LCD_rs_out_w : out std_logic; -- Signal permettant de choisir entre DATA/INSTRUCTION
			LCD_enable_w : out std_logic; -- Signal permettant de valider la commande
			LCD_rw_out_w : out std_logic; -- Signal permettant de s�lectionner le mode write ou read
			LCDD_out_w   : out std_logic_vector(7 downto 0) -- Bus d'instruction vers le LDC
			);
end write_module;


architecture Behavioral of write_module is

	TYPE STATE_TYPE IS (
			READY,
			INIT,
			SIGNAL_SETTLE,
			ENABLE,
			HOLD,
			DONE);

	SIGNAL w_state : STATE_TYPE := READY;
	SIGNAL counter : integer range 0 to 255 := 0; --Compteur d'horloge pour minuter les �tats 100Mhz (T=10 ns)
begin
	process(clk)
	begin

		if rising_edge(clk) then

			case w_state is

				when READY =>
					done_write <= false;

					if (send) then
						w_state <= INIT;
					end if;

				when INIT =>

					-- Pr�pare les signaux qui seront envoy�s au LCD
					LCDD_out_w <= ins_in(7 downto 0);
					LCD_rs_out_w <= ins_in(8);
					LCD_enable_w <= '0';
					LCD_rw_out_w <= '0'; --Mode write

					counter <= 0;

					w_state <= SIGNAL_SETTLE;

				when SIGNAL_SETTLE =>
					LCD_enable_w <= '1';
					w_state <= ENABLE;

				when ENABLE =>

					LCD_enable_w <= '1';

					--Delai d'activation enable 80 ns
					if counter >= 7 then
						w_state <= HOLD;
						counter <= 0;
					else
						counter <= counter + 1;
					end if;

				when HOLD =>

					LCD_enable_w <= '0';

					--Delai avant le prochain write 1200 ns
					if counter >= 119 then
						w_state <= DONE;
						counter <= 0;
					else
						counter <= counter + 1;
					end if;


				when DONE =>

					done_write <= true;

					if (send) then
						w_state <= READY;
					end if;

				when others =>

					w_state <= READY;

			end case;
		end if;
	end process;
end Behavioral;
